`timescale 1ns/1ns
module instmem(input[31:0] address, input clk,rst, output[31:0] inst);
  /*
  reg[31:0] memoryData[0:16383];
 
  
  initial begin
  memoryData[0] = 32'b000000_00001_00010_00000_00000000000;
  memoryData[1] = 32'b000000_00011_00100_00000_00000000000;
  memoryData[2] = 32'b000000_00101_00110_00000_00000000000;
  memoryData[3] = 32'b000000_00111_01000_00010_00000000000;
  memoryData[4] = 32'b000000_01001_01010_00011_00000000000;
  memoryData[5] = 32'b000000_01011_01100_00000_00000000000;
  memoryData[6] = 32'b000000_01101_01110_00000_00000000000;
  end
  assign inst = memoryData[address >> 2];
 */
  logic [31:0] pc, instruction;
  assign pc = address ;
  always@(*) begin
  case (pc)
      0 : instruction <= 32'b11100011101000000000000000010100;
      4 : instruction <= 32'b11100011101000000001101000000001;
      8 : instruction <= 32'b11100011101000000010000100000011;
     12 : instruction <= 32'b11100000100100100011000000000010;
     16 : instruction <= 32'b11100000101000000100000000000000;
     20 : instruction <= 32'b11100000010001000101000100000100;
     24 : instruction <= 32'b11100000110000000110000010100000;
     28 : instruction <= 32'b11100001100001010111000101000010;
     32 : instruction <= 32'b11100000000001111000000000000011;
     36 : instruction <= 32'b11100001111000001001000000000110;
     40 : instruction <= 32'b11100000001001001010000000000101;
     44 : instruction <= 32'b11100001010110000000000000000110;
     48 : instruction <= 32'b00010000100000010001000000000001;
     52 : instruction <= 32'b11100001000110010000000000001000;
     56 : instruction <= 32'b00000000100000100010000000000010;
     60 : instruction <= 32'b11100011101000000000101100000001;
     64 : instruction <= 32'b11100100100000000001000000000000;
     68 : instruction <= 32'b11100100100100001011000000000000; //18
     72 : instruction <= 32'b11100100100000000010000000000100;
     76 : instruction <= 32'b11100100100000000011000000001000;
     80 : instruction <= 32'b11100100100000000100000000001101;
     84 : instruction <= 32'b11100100100000000101000000010000; //22
     88 : instruction <= 32'b11100100100000000110000000010100;
     92 : instruction <= 32'b11100100100100001010000000000100;
     96 : instruction <= 32'b11100100100000000111000000011000; 
    100 : instruction <= 32'b11100011101000000001000000000100; //26 
    104 : instruction <= 32'b11100011101000000010000000000000;
    108 : instruction <= 32'b11100011101000000011000000000000;
    112 : instruction <= 32'b11100000100000000100000100000011; //29
    116 : instruction <= 32'b11100100100101000101000000000000;
    120 : instruction <= 32'b11100100100101000110000000000100;
    124 : instruction <= 32'b11100001010101010000000000000110;
    128 : instruction <= 32'b11000100100001000110000000000000; //33
    132 : instruction <= 32'b11000100100001000101000000000100;
    136 : instruction <= 32'b11100010100000110011000000000001;
    140 : instruction <= 32'b11100011010100110000000000000011; //36
    144 : instruction <= 32'b10111010111111111111111111110111;
    148 : instruction <= 32'b11100010100000100010000000000001;
    152 : instruction <= 32'b11100001010100100000000000000001;
    156 : instruction <= 32'b10111010111111111111111111110011; //40
    160 : instruction <= 32'b11100100100100000001000000000000;
    164 : instruction <= 32'b11100100100100000010000000000100;
    168 : instruction <= 32'b11100100100100000011000000001000; //43
    172 : instruction <= 32'b11100100100100000100000000001100; //44
    176 : instruction <= 32'b11100100100100000101000000010000;
    180 : instruction <= 32'b11100100100100000110000000010100; 
    184 : instruction <= 32'b11101010111111111111111111111111; //47
    default : instruction <= 32'b0; 
  endcase
  end
 assign inst = instruction; 
 
endmodule