`timescale 1ns/1ns

module b32adder(input [31:0] a,b, output reg [31:0] out);
    assign out = a+ b;
endmodule




